magic
tech sky130A
magscale 1 2
timestamp 1641587603
<< nwell >>
rect 1366 442 2276 1080
<< pwell >>
rect 1366 -178 1892 442
<< nmos >>
rect 1566 32 1596 232
rect 1662 32 1692 232
<< pmos >>
rect 1566 661 1596 861
rect 1662 661 1692 861
rect 1758 661 1788 861
rect 1854 661 1884 861
rect 1950 661 1980 861
rect 2046 661 2076 861
<< ndiff >>
rect 1504 220 1566 232
rect 1504 44 1516 220
rect 1550 44 1566 220
rect 1504 32 1566 44
rect 1596 220 1662 232
rect 1596 44 1612 220
rect 1646 44 1662 220
rect 1596 32 1662 44
rect 1692 220 1754 232
rect 1692 44 1708 220
rect 1742 44 1754 220
rect 1692 32 1754 44
<< pdiff >>
rect 1504 849 1566 861
rect 1504 673 1516 849
rect 1550 673 1566 849
rect 1504 661 1566 673
rect 1596 849 1662 861
rect 1596 673 1612 849
rect 1646 673 1662 849
rect 1596 661 1662 673
rect 1692 849 1758 861
rect 1692 673 1708 849
rect 1742 673 1758 849
rect 1692 661 1758 673
rect 1788 849 1854 861
rect 1788 673 1804 849
rect 1838 673 1854 849
rect 1788 661 1854 673
rect 1884 849 1950 861
rect 1884 673 1900 849
rect 1934 673 1950 849
rect 1884 661 1950 673
rect 1980 849 2046 861
rect 1980 673 1996 849
rect 2030 673 2046 849
rect 1980 661 2046 673
rect 2076 849 2138 861
rect 2076 673 2092 849
rect 2126 673 2138 849
rect 2076 661 2138 673
<< ndiffc >>
rect 1516 44 1550 220
rect 1612 44 1646 220
rect 1708 44 1742 220
<< pdiffc >>
rect 1516 673 1550 849
rect 1612 673 1646 849
rect 1708 673 1742 849
rect 1804 673 1838 849
rect 1900 673 1934 849
rect 1996 673 2030 849
rect 2092 673 2126 849
<< psubdiff >>
rect 1402 372 1498 406
rect 1760 372 1856 406
rect 1402 310 1436 372
rect 1822 310 1856 372
rect 1402 -108 1436 -46
rect 1822 -108 1856 -46
rect 1402 -142 1498 -108
rect 1760 -142 1856 -108
<< nsubdiff >>
rect 1402 1010 1498 1044
rect 2144 1010 2240 1044
rect 1402 948 1436 1010
rect 2206 948 2240 1010
rect 1402 512 1436 574
rect 2206 512 2240 574
rect 1402 478 1498 512
rect 2144 478 2240 512
<< psubdiffcont >>
rect 1498 372 1760 406
rect 1402 -46 1436 310
rect 1822 -46 1856 310
rect 1498 -142 1760 -108
<< nsubdiffcont >>
rect 1498 1010 2144 1044
rect 1402 574 1436 948
rect 2206 574 2240 948
rect 1498 478 2144 512
<< poly >>
rect 1566 886 2076 916
rect 1566 861 1596 886
rect 1662 861 1692 886
rect 1758 861 1788 886
rect 1854 861 1884 886
rect 1950 861 1980 886
rect 2046 861 2076 886
rect 1566 636 1596 661
rect 1662 636 1692 661
rect 1758 636 1788 661
rect 1854 636 1884 661
rect 1950 636 1980 661
rect 2046 636 2076 661
rect 1566 630 2076 636
rect 1548 614 2076 630
rect 1548 580 1564 614
rect 1598 606 1756 614
rect 1598 580 1614 606
rect 1548 564 1614 580
rect 1740 580 1756 606
rect 1790 606 1948 614
rect 1790 580 1806 606
rect 1740 564 1806 580
rect 1932 580 1948 606
rect 1982 606 2076 614
rect 1982 580 1998 606
rect 1932 564 1998 580
rect 1644 304 1710 320
rect 1644 284 1660 304
rect 1566 270 1660 284
rect 1694 270 1710 304
rect 1566 254 1710 270
rect 1566 232 1596 254
rect 1662 232 1692 254
rect 1566 10 1596 32
rect 1662 10 1692 32
rect 1566 -20 1692 10
<< polycont >>
rect 1564 580 1598 614
rect 1756 580 1790 614
rect 1948 580 1982 614
rect 1660 270 1694 304
<< locali >>
rect 1402 1010 1498 1044
rect 2144 1010 2240 1044
rect 1402 948 1436 1010
rect 1516 849 1550 865
rect 1516 657 1550 673
rect 1612 849 1646 1010
rect 1612 657 1646 673
rect 1708 849 1742 865
rect 1708 657 1742 673
rect 1804 849 1838 1010
rect 1804 657 1838 673
rect 1900 849 1934 865
rect 1900 657 1934 673
rect 1996 849 2030 1010
rect 2206 948 2240 1010
rect 1996 657 2030 673
rect 2092 849 2126 865
rect 2092 657 2126 673
rect 1548 580 1564 614
rect 1598 580 1614 614
rect 1740 580 1756 614
rect 1790 580 1806 614
rect 1932 580 1948 614
rect 1982 580 1998 614
rect 1402 512 1436 574
rect 2206 512 2240 574
rect 1402 478 1498 512
rect 2144 478 2240 512
rect 1402 372 1498 406
rect 1760 372 1856 406
rect 1402 310 1436 372
rect 1822 310 1856 372
rect 1644 270 1660 304
rect 1694 270 1710 304
rect 1516 220 1550 236
rect 1516 28 1550 44
rect 1612 220 1646 236
rect 1402 -108 1436 -46
rect 1612 -108 1646 44
rect 1708 220 1742 236
rect 1708 28 1742 44
rect 1822 -108 1856 -46
rect 1402 -142 1498 -108
rect 1760 -142 1856 -108
<< viali >>
rect 1516 673 1550 849
rect 1708 673 1742 849
rect 1900 673 1934 849
rect 2092 673 2126 849
rect 1564 580 1598 614
rect 1756 580 1790 614
rect 1948 580 1982 614
rect 1660 270 1694 304
rect 1516 44 1550 220
rect 1708 44 1742 220
<< metal1 >>
rect 1516 861 2126 876
rect 1510 849 2132 861
rect 1510 673 1516 849
rect 1550 848 1708 849
rect 1550 673 1556 848
rect 1510 661 1556 673
rect 1702 673 1708 848
rect 1742 848 1900 849
rect 1742 673 1748 848
rect 1702 661 1748 673
rect 1894 673 1900 848
rect 1934 848 2092 849
rect 1934 673 1940 848
rect 1894 661 1940 673
rect 2086 673 2092 848
rect 2126 673 2132 849
rect 1552 614 1994 620
rect 1552 580 1564 614
rect 1598 580 1756 614
rect 1790 580 1948 614
rect 1982 580 1994 614
rect 1552 574 1994 580
rect 1660 310 1694 574
rect 2086 512 2132 673
rect 1822 478 2132 512
rect 1648 304 1706 310
rect 1648 270 1660 304
rect 1694 270 1706 304
rect 1648 264 1706 270
rect 1510 220 1556 232
rect 1510 44 1516 220
rect 1550 44 1556 220
rect 1702 220 1748 232
rect 1702 44 1708 220
rect 1742 44 1748 220
rect 1822 44 1856 478
rect 1510 32 1856 44
rect 1516 14 1856 32
<< labels >>
rlabel metal1 1674 432 1674 432 7 VIN
port 1 w
rlabel metal1 1838 430 1838 430 7 VOUT
port 2 w
rlabel locali 2224 1024 2224 1024 7 VDD
port 3 w
rlabel locali 1838 -122 1838 -122 7 VSS
port 4 w
<< end >>
