magic
tech sky130A
timestamp 1641260958
<< nwell >>
rect 683 221 1138 540
<< pwell >>
rect 683 -89 946 221
<< nmos >>
rect 783 16 798 116
rect 831 16 846 116
<< pmos >>
rect 783 331 798 431
rect 831 331 846 431
rect 879 331 894 431
rect 927 331 942 431
rect 975 331 990 431
rect 1023 331 1038 431
<< ndiff >>
rect 752 110 783 116
rect 752 22 758 110
rect 775 22 783 110
rect 752 16 783 22
rect 798 110 831 116
rect 798 22 806 110
rect 823 22 831 110
rect 798 16 831 22
rect 846 110 877 116
rect 846 22 854 110
rect 871 22 877 110
rect 846 16 877 22
<< pdiff >>
rect 752 424 783 431
rect 752 336 758 424
rect 775 336 783 424
rect 752 331 783 336
rect 798 424 831 431
rect 798 336 806 424
rect 823 336 831 424
rect 798 331 831 336
rect 846 424 879 431
rect 846 336 854 424
rect 871 336 879 424
rect 846 331 879 336
rect 894 424 927 431
rect 894 336 902 424
rect 919 336 927 424
rect 894 331 927 336
rect 942 424 975 431
rect 942 336 950 424
rect 967 336 975 424
rect 942 331 975 336
rect 990 424 1023 431
rect 990 336 998 424
rect 1015 336 1023 424
rect 990 331 1023 336
rect 1038 424 1069 431
rect 1038 336 1046 424
rect 1063 336 1069 424
rect 1038 331 1069 336
<< ndiffc >>
rect 758 22 775 110
rect 806 22 823 110
rect 854 22 871 110
<< pdiffc >>
rect 758 336 775 424
rect 806 336 823 424
rect 854 336 871 424
rect 902 336 919 424
rect 950 336 967 424
rect 998 336 1015 424
rect 1046 336 1063 424
<< psubdiff >>
rect 701 186 749 203
rect 880 186 928 203
rect 701 155 718 186
rect 911 155 928 186
rect 701 -54 718 -23
rect 911 -54 928 -23
rect 701 -71 749 -54
rect 880 -71 928 -54
<< nsubdiff >>
rect 701 505 749 522
rect 1072 505 1120 522
rect 701 474 718 505
rect 1103 474 1120 505
rect 701 256 718 287
rect 1103 256 1120 287
rect 701 239 749 256
rect 1072 239 1120 256
<< psubdiffcont >>
rect 749 186 880 203
rect 701 -23 718 155
rect 911 -23 928 155
rect 749 -71 880 -54
<< nsubdiffcont >>
rect 749 505 1072 522
rect 701 287 718 474
rect 1103 287 1120 474
rect 749 239 1072 256
<< poly >>
rect 783 443 1038 458
rect 783 431 798 443
rect 831 431 846 443
rect 879 431 894 443
rect 927 431 942 443
rect 975 431 990 443
rect 1023 431 1038 443
rect 783 318 798 331
rect 831 318 846 331
rect 879 318 894 331
rect 927 318 942 331
rect 975 318 990 331
rect 1023 318 1038 331
rect 783 315 1038 318
rect 774 307 1038 315
rect 774 290 782 307
rect 799 303 878 307
rect 799 290 807 303
rect 774 282 807 290
rect 870 290 878 303
rect 895 303 974 307
rect 895 290 903 303
rect 870 282 903 290
rect 966 290 974 303
rect 991 303 1038 307
rect 991 290 999 303
rect 966 282 999 290
rect 822 152 855 160
rect 822 142 830 152
rect 783 135 830 142
rect 847 135 855 152
rect 783 127 855 135
rect 783 116 798 127
rect 831 116 846 127
rect 783 5 798 16
rect 831 5 846 16
rect 783 -10 846 5
<< polycont >>
rect 782 290 799 307
rect 878 290 895 307
rect 974 290 991 307
rect 830 135 847 152
<< locali >>
rect 701 505 749 522
rect 1072 505 1120 522
rect 701 474 718 505
rect 746 480 775 488
rect 763 463 775 480
rect 758 424 775 463
rect 758 328 775 336
rect 806 480 823 488
rect 823 463 1015 475
rect 806 458 1015 463
rect 806 424 823 458
rect 806 328 823 336
rect 854 424 871 432
rect 854 328 871 336
rect 902 424 919 458
rect 902 328 919 336
rect 950 424 967 432
rect 950 328 967 336
rect 998 424 1015 458
rect 1103 474 1120 505
rect 998 328 1015 336
rect 1046 424 1063 432
rect 1046 328 1063 336
rect 774 290 782 307
rect 799 290 807 307
rect 870 290 878 307
rect 895 290 903 307
rect 966 290 974 307
rect 991 290 999 307
rect 701 256 718 287
rect 1120 287 1163 336
rect 1103 256 1163 287
rect 701 239 749 256
rect 1072 246 1163 256
rect 1072 239 1120 246
rect 701 186 749 203
rect 880 186 928 203
rect 701 155 718 186
rect 911 181 928 186
rect 911 155 1163 181
rect 822 135 830 152
rect 847 135 855 152
rect 758 110 775 118
rect 758 -11 775 22
rect 701 -54 718 -23
rect 746 -19 775 -11
rect 763 -36 775 -19
rect 806 110 823 118
rect 806 -19 823 22
rect 854 110 871 118
rect 854 14 871 22
rect 928 91 1163 155
rect 1353 67 1380 71
rect 1353 50 1357 67
rect 1374 50 1380 67
rect 1353 46 1380 50
rect 911 -54 928 -23
rect 701 -71 749 -54
rect 880 -71 928 -54
<< viali >>
rect 746 463 763 480
rect 758 336 775 424
rect 806 463 823 480
rect 854 336 871 424
rect 950 336 967 424
rect 1046 336 1063 424
rect 782 290 799 307
rect 878 290 895 307
rect 974 290 991 307
rect 830 135 847 152
rect 758 22 775 110
rect 746 -36 763 -19
rect 854 22 871 110
rect 806 -36 823 -19
rect 1142 50 1159 67
rect 1357 50 1374 67
<< metal1 >>
rect 738 485 771 488
rect 738 458 741 485
rect 768 458 771 485
rect 738 455 771 458
rect 798 485 831 488
rect 798 458 801 485
rect 828 458 831 485
rect 798 455 831 458
rect 758 430 1063 438
rect 755 424 1066 430
rect 755 336 758 424
rect 775 336 778 424
rect 755 330 778 336
rect 851 336 854 424
rect 871 336 874 424
rect 851 330 874 336
rect 947 336 950 424
rect 967 336 970 424
rect 947 330 970 336
rect 1043 336 1046 424
rect 1063 336 1066 424
rect 1043 330 1066 336
rect 776 307 1026 310
rect 776 290 782 307
rect 799 290 878 307
rect 895 290 974 307
rect 991 290 1026 307
rect 776 287 1026 290
rect 997 226 1026 287
rect 997 197 1441 226
rect 822 152 1055 160
rect 822 135 830 152
rect 847 135 1055 152
rect 822 131 1055 135
rect 755 110 778 116
rect 755 22 758 110
rect 775 22 778 110
rect 851 110 874 116
rect 851 22 854 110
rect 871 22 874 110
rect 1026 73 1055 131
rect 1412 73 1441 197
rect 1026 67 1165 73
rect 1026 50 1142 67
rect 1159 50 1165 67
rect 1026 44 1165 50
rect 1351 67 1441 73
rect 1351 50 1357 67
rect 1374 50 1441 67
rect 1351 43 1441 50
rect 755 16 896 22
rect 758 7 896 16
rect 738 -14 771 -11
rect 738 -41 741 -14
rect 768 -41 771 -14
rect 738 -44 771 -41
rect 798 -14 831 -11
rect 798 -41 801 -14
rect 828 -41 831 -14
rect 798 -44 831 -41
<< via1 >>
rect 741 480 768 485
rect 741 463 746 480
rect 746 463 763 480
rect 763 463 768 480
rect 741 458 768 463
rect 801 480 828 485
rect 801 463 806 480
rect 806 463 823 480
rect 823 463 828 480
rect 801 458 828 463
rect 741 -19 768 -14
rect 741 -36 746 -19
rect 746 -36 763 -19
rect 763 -36 768 -19
rect 741 -41 768 -36
rect 801 -19 828 -14
rect 801 -36 806 -19
rect 806 -36 823 -19
rect 823 -36 828 -19
rect 801 -41 828 -36
<< metal2 >>
rect 738 485 772 488
rect 738 458 741 485
rect 768 458 772 485
rect 738 -14 772 458
rect 738 -41 741 -14
rect 768 -41 772 -14
rect 738 -44 772 -41
rect 798 485 831 488
rect 798 458 801 485
rect 828 458 831 485
rect 798 -14 831 458
rect 798 -41 801 -14
rect 828 -41 831 -14
rect 798 -44 831 -41
use INVMIN_v1p1  INVMIN_v1p1_0
timestamp 1641260958
transform 1 0 1288 0 1 96
box -150 -75 85 265
<< labels >>
flabel via1 754 470 754 470 0 FreeSans 240 0 0 0 VIN
port 0 nsew
flabel via1 816 -27 816 -27 0 FreeSans 240 0 0 0 VOUT
port 1 nsew
flabel metal1 883 144 883 144 0 FreeSans 240 0 0 0 CTR
port 2 nsew
flabel locali 1148 294 1148 294 0 FreeSans 240 0 0 0 VDD
port 3 nsew
flabel locali 1103 136 1103 136 0 FreeSans 240 0 0 0 VSS
port 4 nsew
<< end >>
