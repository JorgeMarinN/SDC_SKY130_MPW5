magic
tech sky130A
magscale 1 2
timestamp 1640034244
<< error_p >>
rect -173 181 -115 187
rect 19 181 77 187
rect 211 181 269 187
rect -173 147 -161 181
rect 19 147 31 181
rect 211 147 223 181
rect -173 141 -115 147
rect 19 141 77 147
rect 211 141 269 147
rect -269 -147 -211 -141
rect -77 -147 -19 -141
rect 115 -147 173 -141
rect -269 -181 -257 -147
rect -77 -181 -65 -147
rect 115 -181 127 -147
rect -269 -187 -211 -181
rect -77 -187 -19 -181
rect 115 -187 173 -181
<< nwell >>
rect -455 -319 455 319
<< pmos >>
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
<< pdiff >>
rect -317 88 -255 100
rect -317 -88 -305 88
rect -271 -88 -255 88
rect -317 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 317 100
rect 255 -88 271 88
rect 305 -88 317 88
rect 255 -100 317 -88
<< pdiffc >>
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
<< nsubdiff >>
rect -419 249 -323 283
rect 323 249 419 283
rect -419 187 -385 249
rect 385 187 419 249
rect -419 -249 -385 -187
rect 385 -249 419 -187
rect -419 -283 -323 -249
rect 323 -283 419 -249
<< nsubdiffcont >>
rect -323 249 323 283
rect -419 -187 -385 187
rect 385 -187 419 187
rect -323 -283 323 -249
<< poly >>
rect -177 181 -111 197
rect -177 147 -161 181
rect -127 147 -111 181
rect -177 131 -111 147
rect 15 181 81 197
rect 15 147 31 181
rect 65 147 81 181
rect 15 131 81 147
rect 207 181 273 197
rect 207 147 223 181
rect 257 147 273 181
rect 207 131 273 147
rect -255 100 -225 126
rect -159 100 -129 131
rect -63 100 -33 126
rect 33 100 63 131
rect 129 100 159 126
rect 225 100 255 131
rect -255 -131 -225 -100
rect -159 -126 -129 -100
rect -63 -131 -33 -100
rect 33 -126 63 -100
rect 129 -131 159 -100
rect 225 -126 255 -100
rect -273 -147 -207 -131
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -273 -197 -207 -181
rect -81 -147 -15 -131
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect -81 -197 -15 -181
rect 111 -147 177 -131
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 111 -197 177 -181
<< polycont >>
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
<< locali >>
rect -419 249 -323 283
rect 323 249 419 283
rect -419 187 -385 249
rect 385 187 419 249
rect -177 147 -161 181
rect -127 147 -111 181
rect 15 147 31 181
rect 65 147 81 181
rect 207 147 223 181
rect 257 147 273 181
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect 111 -181 127 -147
rect 161 -181 177 -147
rect -419 -249 -385 -187
rect 385 -249 419 -187
rect -419 -283 -323 -249
rect 323 -283 419 -249
<< viali >>
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
<< metal1 >>
rect -173 181 -115 187
rect -173 147 -161 181
rect -127 147 -115 181
rect -173 141 -115 147
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect 211 181 269 187
rect 211 147 223 181
rect 257 147 269 181
rect 211 141 269 147
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect -269 -147 -211 -141
rect -269 -181 -257 -147
rect -223 -181 -211 -147
rect -269 -187 -211 -181
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -31 -181 -19 -147
rect -77 -187 -19 -181
rect 115 -147 173 -141
rect 115 -181 127 -147
rect 161 -181 173 -147
rect 115 -187 173 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -402 -266 402 266
string parameters w 1 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
