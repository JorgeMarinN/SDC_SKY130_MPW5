magic
tech sky130A
timestamp 1641587603
<< locali >>
rect 9731 2964 9837 3014
rect 9731 2911 9741 2964
rect 9827 2911 9837 2964
rect 10152 2991 10264 3014
rect 10152 2938 10165 2991
rect 10251 2938 10264 2991
rect 10152 2923 10264 2938
rect 9731 2901 9837 2911
<< viali >>
rect 9741 2911 9827 2964
rect 10165 2938 10251 2991
<< metal1 >>
rect 9556 3243 9732 3279
rect 2500 3187 9732 3243
rect 9556 3186 9732 3187
rect 9732 3023 10202 3034
rect 9732 3022 10046 3023
rect 9731 2964 9837 2975
rect 9731 2911 9741 2964
rect 9827 2911 9837 2964
rect 9731 2901 9837 2911
rect 9888 2635 10046 3022
rect 10152 2991 10264 3000
rect 10152 2938 10165 2991
rect 10251 2938 10264 2991
rect 10152 2923 10264 2938
rect 9888 2634 10202 2635
rect 2361 2584 10478 2634
<< via1 >>
rect 9741 2911 9827 2964
rect 10165 2938 10251 2991
<< metal2 >>
rect 1982 3296 9647 3380
rect 1982 2754 2066 3296
rect 2563 2752 5566 2838
rect 6063 2752 9066 2838
rect 9563 2752 9647 3296
rect 10152 2991 10264 3000
rect 9731 2964 9837 2975
rect 9731 2911 9741 2964
rect 9827 2911 9837 2964
rect 10152 2938 10165 2991
rect 10251 2938 10264 2991
rect 10152 2923 10264 2938
rect 9731 2901 9837 2911
rect 8980 2681 9066 2752
rect 9751 2681 9837 2901
rect 8979 2595 9838 2681
<< metal3 >>
rect 1420 2501 1500 2581
rect 4920 2501 5000 2581
rect 8420 2501 8500 2581
<< metal5 >>
rect 196 2791 2928 2951
rect 3696 2791 6428 2951
rect 7196 2791 9468 2951
use BUFFMIN_v1p1  BUFFMIN_v1p1_0
timestamp 1641587603
transform 1 0 9747 0 1 2969
box -15 -5 455 335
use INVandCAP_v1p1  INVandCAP_v1p1_2
timestamp 1641587603
transform 1 0 6994 0 1 5
box 0 0 3484 3238
use INVandCAP_v1p1  INVandCAP_v1p1_1
timestamp 1641587603
transform 1 0 3494 0 1 5
box 0 0 3484 3238
use INVandCAP_v1p1  INVandCAP_v1p1_0
timestamp 1641587603
transform 1 0 -6 0 1 5
box 0 0 3484 3238
<< labels >>
flabel metal1 2813 3212 2813 3212 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal1 2756 2602 2756 2602 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal2 2024 3333 2024 3333 0 FreeSans 800 0 0 0 SENS_IN
port 3 nsew
flabel metal2 3520 2790 3520 2790 0 FreeSans 800 0 0 0 N1
port 4 nsew
flabel metal5 8006 2877 8006 2877 0 FreeSans 800 0 0 0 CON_CV
port 6 nsew
flabel locali 10181 3000 10181 3000 0 FreeSans 800 0 0 0 N2
port 7 nsew
<< end >>
