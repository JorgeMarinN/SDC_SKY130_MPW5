magic
tech sky130A
magscale 1 2
timestamp 1640196996
<< metal4 >>
rect -2399 2279 2399 2320
rect -2399 -2279 2143 2279
rect 2379 -2279 2399 2279
rect -2399 -2320 2399 -2279
<< via4 >>
rect 2143 -2279 2379 2279
<< mimcap2 >>
rect -2299 2180 2141 2220
rect -2299 -2180 -239 2180
rect 81 -2180 2141 2180
rect -2299 -2220 2141 -2180
<< mimcap2contact >>
rect -239 -2180 81 2180
<< metal5 >>
rect 2101 2279 2421 2321
rect -263 2180 105 2204
rect -263 -2180 -239 2180
rect 81 -2180 105 2180
rect -263 -2204 105 -2180
rect 2101 -2279 2143 2279
rect 2379 -2279 2421 2279
rect 2101 -2321 2421 -2279
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2399 -2320 2241 2320
string parameters w 22.2 l 22.2 val 1.002k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 5
string library sky130
<< end >>
