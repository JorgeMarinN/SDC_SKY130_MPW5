magic
tech sky130A
magscale 1 2
timestamp 1641588824
<< nwell >>
rect 20800 8076 20998 8234
rect 20734 7666 21644 8076
<< locali >>
rect 22756 7244 22816 7260
<< viali >>
rect 20866 7630 21512 7664
rect 22756 7260 22816 7320
rect 21874 6568 21934 6628
rect 21224 6444 21284 6504
<< metal1 >>
rect 7826 9164 7920 9222
rect 22668 9130 23616 9242
rect 7778 7942 7862 7996
rect 20866 7676 21514 7848
rect 22122 7806 22774 8026
rect 23558 7818 23616 9130
rect 22788 7750 22864 7766
rect 22788 7698 22795 7750
rect 22847 7698 22864 7750
rect 22788 7692 22864 7698
rect 20858 7664 21522 7676
rect 20858 7630 20866 7664
rect 21512 7630 21522 7664
rect 20858 7616 21522 7630
rect 23558 7658 23638 7818
rect 23558 7600 23616 7658
rect 23558 7564 23638 7600
rect 22744 7320 22828 7332
rect 22744 7260 22756 7320
rect 22816 7260 22828 7320
rect 22744 7248 22828 7260
rect 21862 6628 21946 6640
rect 21862 6568 21874 6628
rect 21934 6568 21946 6628
rect 21862 6556 21946 6568
rect 21212 6504 21298 6518
rect 21212 6444 21224 6504
rect 21284 6444 21298 6504
rect 21212 6430 21298 6444
rect 23528 6408 23616 6444
rect 23528 6248 23638 6408
rect 22590 6224 23094 6232
rect 22122 6004 23094 6224
rect 23528 5874 23616 6248
rect 22106 5864 23616 5874
rect 22106 5804 22182 5864
rect 22242 5804 23616 5864
rect 22106 5794 23616 5804
<< via1 >>
rect 22795 7698 22847 7750
rect 22756 7260 22816 7320
rect 21874 6568 21934 6628
rect 21224 6444 21284 6504
rect 22182 5804 22242 5864
<< metal2 >>
rect 9142 7660 9374 7780
rect 22022 7756 22246 8434
rect 22022 7750 22854 7756
rect 22022 7698 22795 7750
rect 22847 7698 22854 7750
rect 22022 7692 22854 7698
rect 20790 7562 20912 7644
rect 20998 7514 21102 7562
rect 20998 7056 21006 7514
rect 21092 7056 21102 7514
rect 20998 7046 21102 7056
rect 22402 7320 22822 7328
rect 22402 7260 22756 7320
rect 22816 7260 22822 7320
rect 22402 7254 22822 7260
rect 22402 6636 22476 7254
rect 21868 6628 22476 6636
rect 21868 6568 21874 6628
rect 21934 6568 22476 6628
rect 21868 6562 22476 6568
rect 21218 6504 22248 6510
rect 21218 6444 21224 6504
rect 21284 6444 22248 6504
rect 21218 6438 22248 6444
rect 22176 5864 22248 6438
rect 22176 5804 22182 5864
rect 22242 5804 22248 5864
rect 22176 5798 22248 5804
rect 22994 5626 23062 6528
rect 22220 5472 23062 5626
<< via2 >>
rect 21006 7056 21092 7514
<< metal3 >>
rect 20998 7514 21102 7562
rect 20998 7056 21006 7514
rect 21092 7056 21102 7514
rect 20998 7046 21102 7056
<< via3 >>
rect 21006 7056 21092 7514
<< metal4 >>
rect 20620 8356 21102 8502
rect 20420 8320 21102 8356
rect 20998 7514 21102 8320
rect 20998 7056 21006 7514
rect 21092 7056 21102 7514
rect 20998 7046 21102 7056
<< via4 >>
rect 20384 8356 20620 8592
<< metal5 >>
rect 20280 8592 20514 8676
rect 20280 8356 20384 8592
rect 20620 8356 20654 8504
rect 20280 8320 20654 8356
rect 20654 5208 21574 5528
use DFF_v4p1  DFF_v4p1_0
timestamp 1641579593
transform 0 -1 23156 1 0 6824
box -636 -618 1036 626
use PASSGATE_v1p2  PASSGATE_v1p2_0
timestamp 1641260958
transform 1 0 19368 0 1 6586
box 1366 -178 2882 1080
use OSC_v3p2  OSC_v3p2_1
timestamp 1641587603
transform 1 0 1718 0 -1 14404
box -12 10 20956 6760
use OSC_v3p2  OSC_v3p2_0
timestamp 1641587603
transform 1 0 1718 0 1 -374
box -12 10 20956 6760
<< labels >>
flabel metal1 7808 7968 7808 7968 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 7874 9190 7874 9190 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal2 9244 7732 9244 7732 0 FreeSans 1600 0 0 0 SENS_IN
port 2 nsew
flabel metal5 20956 5398 20956 5398 0 FreeSans 1600 0 0 0 REF_IN
port 3 nsew
flabel metal2 22458 7288 22458 7288 0 FreeSans 1600 0 0 0 DOUT
port 4 nsew
<< end >>
