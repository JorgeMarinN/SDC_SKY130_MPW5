magic
tech sky130A
magscale 1 2
timestamp 1640649115
<< metal3 >>
rect -2016 2292 2016 2320
rect -2016 -2292 1932 2292
rect 1996 -2292 2016 2292
rect -2016 -2320 2016 -2292
<< via3 >>
rect 1932 -2292 1996 2292
<< mimcap >>
rect -1916 2180 1844 2220
rect -1916 -2180 -128 2180
rect 56 -2180 1844 2180
rect -1916 -2220 1844 -2180
<< mimcapcontact >>
rect -128 -2180 56 2180
<< metal4 >>
rect 1916 2292 2012 2308
rect -129 2180 57 2181
rect -129 -2180 -128 2180
rect 56 -2180 57 2180
rect -129 -2181 57 -2180
rect 1916 -2292 1932 2292
rect 1996 -2292 2012 2292
rect 1916 -2308 2012 -2292
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -2016 -2320 1944 2320
string parameters w 18.8 l 22.2 val 850.3 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 5
string library sky130
<< end >>
