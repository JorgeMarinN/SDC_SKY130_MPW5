magic
tech sky130A
magscale 1 2
timestamp 1641587603
<< error_s >>
rect 6000 4640 6080 4720
rect 5920 4560 6000 4640
<< metal2 >>
rect 9938 4612 10022 4622
rect 9938 28 9948 4612
rect 10012 28 10022 4612
rect 9938 18 10022 28
<< via2 >>
rect 9948 28 10012 4612
<< metal3 >>
rect 6000 5160 6320 5190
rect 6000 4924 6042 5160
rect 6278 4924 6320 5160
rect 6000 4640 6320 4924
rect 5016 4612 10032 4640
rect 5016 4374 9948 4612
rect 6000 28 9948 4374
rect 10012 28 10032 4612
rect 4130 -110 4414 2
rect 6000 0 10032 28
rect 4130 -346 4156 -110
rect 4392 -346 4414 -110
rect 4130 -432 4414 -346
<< via3 >>
rect 6042 4924 6278 5160
rect 4156 -346 4392 -110
<< mimcap >>
rect 6100 4500 9860 4540
rect 6100 140 9636 4500
rect 9820 140 9860 4500
rect 6100 100 9860 140
<< mimcapcontact >>
rect 9636 140 9820 4500
<< metal4 >>
rect 8628 5268 9822 5306
rect 6000 5160 6320 5190
rect 3470 5094 4558 5142
rect 3470 4858 3506 5094
rect 3742 4858 4558 5094
rect 3470 4826 4558 4858
rect 4490 4498 4558 4826
rect 6000 4924 6042 5160
rect 6278 4924 6320 5160
rect 8848 5014 9822 5268
rect 6000 4640 6320 4924
rect 9634 4500 9822 5014
rect 9634 140 9636 4500
rect 9820 140 9822 4500
rect 9634 138 9822 140
rect 4130 -110 4414 2
rect 4130 -346 4156 -110
rect 4392 -346 4414 -110
rect 4130 -432 4414 -346
<< via4 >>
rect 3506 4858 3742 5094
rect 8612 5032 8848 5268
<< metal5 >>
rect 8526 5268 8936 5306
rect 3472 5094 3792 5140
rect 3472 4858 3506 5094
rect 3742 4858 3792 5094
rect 3472 4524 3792 4858
rect 8526 5032 8612 5268
rect 8848 5032 8936 5268
rect 3472 4500 3506 4524
rect 8526 4500 8936 5032
use sky130_fd_pr__cap_mim_m3_2_7PBNAZ  sky130_fd_pr__cap_mim_m3_2_7PBNAZ_0
timestamp 1640651334
transform 1 0 3739 0 1 2320
box -671 -2321 693 2321
use sky130_fd_pr__cap_mim_m3_1_9K4XRG  sky130_fd_pr__cap_mim_m3_1_9K4XRG_0
timestamp 1640651334
transform 1 0 4560 0 1 2320
box -456 -2320 456 2320
use sky130_fd_pr__cap_mim_m3_2_4SGG6N  sky130_fd_pr__cap_mim_m3_2_4SGG6N_0
timestamp 1641587603
transform 1 0 7323 0 1 2320
box -2231 -2321 2253 2321
<< labels >>
flabel metal4 6140 4764 6140 4764 0 FreeSans 1600 0 0 0 BOT
port 2 nsew
flabel metal4 9210 5152 9210 5152 0 FreeSans 1600 0 0 0 TOP_B
port 4 nsew
flabel metal4 4110 4986 4110 4986 0 FreeSans 1600 0 0 0 TOP_V
port 3 nsew
<< end >>
